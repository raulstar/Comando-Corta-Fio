* COMANDO CORTA FIO                             Revised: Friday, March 17, 2000
* C:\MEUS DOCUMENTOS\MEUS DOCUMENTOS\COMANDO CORRevision: RAUL
* ELETRONICA RACIONAL
* RUA VITAL BRASIL n02 J. TUP� BARUERI
* 
* 
* 
120V 8581 0 
+12 8586 0 
+5 8593 0 
GND_POWER 8595 0 
Q6 8599 8589 8593 BC548
K2 8581  8585 8586 8582 GUILHOTINA
U1 8599 8596 8591 8594 8592 8597 8598 8591       8593 8595 4017
U2 8586 8580 8593 LM78L05ACZ
R1 8596 8595 1M
R2 8599 8595 1M
R3 8591 8595 1M
R4 8598 8600 100K
R5 8597 8590 100K
R6 8580 8595 470r
R7 8594 8589 100K
R8 8587 8600 100K
R9 8588 8601 100K
C1 8600 8595 1uF
C2 8590 8595 4,7uF
C3 8601 8595 4,7uF
C4 8589 8595 1uF
C5 8593 8595 1000uF
C6 8593 8595 100nf
C7 8586 8595 2200uF
JP1 8595 8599 8591 8596 8593 CONTROLE
JP2 8581 8584 8585 SAIDA
JP3 8595 8578 8579 TRAFO
JP4 8592 8601 AJUSTE
R10 8580 8593 220r
D1 8600 8598 1N4004
D2 8590 8597 1N4004
D3 8601 8592 1N4004
D4 8589 8594 1N4004
D5 8579 8586 1N4004
D6 8578 8586 1N4004
D7 8583 8586 1N4004
D8 8582 8586 1N4004
Q1 8599 8600 8593 BC548
Q2 8595 8587 8582 BC548
Q3 8599 8590 8593 BC548
Q4 8599 8601 8593 BC548
Q5 8595 8588 8583 BC548
K1 8581  8584 8586 8583 MOTOR
.END
